package frontend_pkg;

typedef struct packed {
        logic valid;
        logic taken;
    } bht_prediction_t;

endpackage